module dut();

endmodule
