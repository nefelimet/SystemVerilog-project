module test_dut;


endmodule
